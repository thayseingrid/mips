library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoria_instrucao is
    port (
        endereco  : in std_logic_vector(5 downto 0);
        instrucao : out std_logic_vector(31 downto 0)
    );
end memoria_instrucao;

architecture memoria_instrucao of memoria_instrucao is
    type tipo_ram is array (0 to 63) of std_logic_vector(31 downto 0);

    signal ram : tipo_ram;
begin
    ram <= (
        -- add r1, r0, r0
        0 => "000000" & "00000" & "00000" & "00001" & "00000" & "100000",

        -- add r2, r0, r0
        1 => "000000" & "00000" & "00000" & "00010" & "00000" & "100000",

        -- addi r3, r0, 10
        2 => "001000" & "00000" & "00011" & "0000000000001010",
 
        -- slt r8, r1, r3
        3 => "000000" & "00001" & "00011" & "01000" & "00000" & "101010",

        -- add r0, r0, r0
        4 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",
        
        -- add r0, r0, r0
        5 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0
        6 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- beq r8, r0, fim
        7 => "000100" & "01000" & "00000" & "0000000000010001",
        
        -- add r0, r0, r0
        8 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0      
        9 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0
        10 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r8, r1, r7
        11 => "000000" & "00001" & "00111" & "01000" & "00000" & "100000",

        -- add r0, r0, r0
        12 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0      
        13 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0
        14 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- sw r2, 0(r8)
        15 => "101011" & "01000" & "00010" & "0000000000000000",

        -- addi r1, r1, 1
        16 => "001000" & "00001" & "00001" & "0000000000000001",

        -- add r0, r0, r0
        17 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0      
        18 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0
        19 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r2, r2, r1
        20 => "000000" & "00010" & "00001" & "00010" & "00000" & "100000",

        -- j enquanto
        21 => "000010" & "11111111111111111111101101",

        -- add r0, r0, r0
        22 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0      
        23 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- add r0, r0, r0
        24 => "000000" & "00000" & "00000" & "00000" & "00000" & "100000",

        -- lw r2, 9(r7)
        25 => "100011" & "00111" & "00010" & "0000000000001001",

        
        others => "000000" & "00000" & "00000" & "00000" & "00000" & "100000"
    );


    process (endereco)
    begin
        instrucao <= ram(to_integer(unsigned(endereco))); --instrucao = ram[endereco]
    end process;
end memoria_instrucao;
